module top (
    input wire clk
);

  // instr fetch signals
  wire [31:0] instr;
  wire pc_enable;
  wire pc_load;
  wire [31:0] load_addr;
  wire [31:0] pc_out;

  // control signals from decoder
  wire [3:0] alu_ops;
  wire reg_write;
  wire mem_read;
  wire mem_write;
  wire [1:0] mem_width;
  wire is_branch;
  wire [2:0] branch_type;
  wire is_jump;
  wire is_jalr;
  wire [4:0] rs1;
  wire [4:0] rs2;
  wire rs1_used;
  wire rs2_used;
  wire [4:0] rd;
  wire [31:0] imm;

  // pc control
  assign pc_enable = 1'b1;
  assign pc_load   = 1'b0;  // modify this based on branch/jump results
  assign load_addr = 32'b0;  // set this to branch/jump target

  // reset logic
  reg rst;
  initial begin
    rst = 1'b1;
    #10 rst = 1'b0;
  end

  program_counter pc_inst (
      .clk(clk),
      .rst(rst),
      .enable(pc_enable),
      .load(pc_load),
      .addr(load_addr),
      .pc(pc_out)
  );

  instruction_memory instr_mem (
      .addr(pc_out),
      .instr_out(instr)
  );

  decoder decoder_inst (
      .instr(instr),
      .alu_ops(alu_ops),
      .reg_write(reg_write),
      .mem_read(mem_read),
      .mem_write(mem_write),
      .mem_width(mem_width),
      .is_branch(is_branch),
      .branch_type(branch_type),
      .is_jump(is_jump),
      .is_jalr(is_jalr),
      .rs1(rs1),
      .rs2(rs2),
      .rs1_used(rs1_used),
      .rs2_used(rs2_used),
      .rd(rd),
      .imm(imm)
  );

endmodule
